*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../ciceda/models/ptm_130_ngspice.spi
.include ../../../ciceda/lib/SUN_TR_GF130N.spi
.include ../../../ciceda/lib/SUN_TRIO_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc 1.5
VSS VSS 0 dc 0

V1 ERASE VSS PULSE(0, 1.5, 0, 10n, 10n, 600n, 1200u, 0) dc 0
V2 EXPOSE VSS PULSE(0, 1.5, 600n, 10n, 10n, 30u, 1200u, 0) dc 0
V3 VRESET VSS dc 1.5

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include sensor.cir
XDUT VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------

.control
set color0=white
set color1=black
tran 1n 1200u
plot V(VSTORE) V(EXPOSE) V(ERASE) V(XDUT.VPG)
wrdata ../output/tb_sensor_settle.txt V(VSTORE) V(EXPOSE) V(ERASE) V(XDUT.VPG) @m.xdut.m2[id] @m.xdut.m2[gm]
.endc
.end
