.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

X1 VCMP_OUT DATA_0 READ VSS MEMCELL
X2 VCMP_OUT DATA_1 READ VSS MEMCELL
X3 VCMP_OUT DATA_2 READ VSS MEMCELL
X4 VCMP_OUT DATA_3 READ VSS MEMCELL
X5 VCMP_OUT DATA_4 READ VSS MEMCELL
X6 VCMP_OUT DATA_5 READ VSS MEMCELL
X7 VCMP_OUT DATA_6 READ VSS MEMCELL
X8 VCMP_OUT DATA_7 READ VSS MEMCELL

.ENDS

.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
V1 VS VSS dc 0
.ENDS