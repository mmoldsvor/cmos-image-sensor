.SUBCKT PIXEL_SENSOR VCLK VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

.include sensor.cir
X1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

.include comp_improved_dynamic.cir
X2 VSTORE VRAMP VCLK VOUTP VOUTN VDD VSS COMP

*.include sr_latch.cir
*XSR1 VOUTN VSS Q QN VDD VSS SR

.include memory.cir
X3 READ VSS DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS