*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../ciceda/models/ptm_130_ngspice.spi
.include ../../../ciceda/lib/SUN_TR_GF130N.spi
.include ../../../ciceda/lib/SUN_TRIO_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc 1.5
V1 VSTORE VSS dc 0.7
VSS VSS 0 dc 0
V2 VRAMP VSS PULSE(0, 1.5, 0, 60u, 10n, 60u, 120u, 0) dc 0
V3 VCLK VSS PULSE(0, 1.5, 500n, 1n, 1n, 500n, 1u, 0) dc 0
V4 VRESET VSS PULSE(0, 1.5, 25u, 1n, 1n, 60u, 60u, 0) dc 0

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include comp_improved_dynamic.cir
XDUT VSTORE VRAMP VCLK VOUTP VOUTN VDD VSS COMP

XSR1 VOUTN VCLK VRESET Q QN VDD VSS DFRNQNX1_CV

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------

.control
set color0=white
set color1=black
tran 1n 60u
plot V(VSTORE) V(VRAMP) V(VOUTP) V(VOUTN) V(VCLK)
wrdata ../output/tb_comp.txt V(VSTORE) V(VRAMP) V(VOUTP) V(VOUTN) V(VCLK) V(VRESET) V(Q) V(QN)
.endc
.end
