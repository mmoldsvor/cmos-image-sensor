*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../ciceda/models/ptm_130_ngspice.spi
.include ../../../ciceda/lib/SUN_TR_GF130N.spi
.include ../../../ciceda/lib/SUN_TRIO_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc 1.5
VSS VSS 0 dc 0
V1 IO VSS PULSE(0, 1.5, 0, 10n, 10n, 7.5u, 30u, 0) dc 0
V2 READ VSS PULSE(0, 1.5, 15u, 10n, 10n, 10u, 30u, 0) dc 0
V3 VCMP_OUT VSS PULSE(0, 1.5, 40u, 10n, 10n, 2.5u, 60u, 0) dc 0

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include memory.cir
M1 DATA_0 IO VDD VDD pmos w=0.5u l=0.5u
XDUT VCMP_OUT DATA_0 READ VSS MEMCELL

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------

.control
set color0=white
set color1=black
tran 1n 60u
plot V(VCMP_OUT) V(DATA_0) V(READ) V(XDUT.vg) V(XDUT.dmem)
wrdata ../output/tb_memcell.txt V(VCMP_OUT) V(DATA_0), V(IO) V(READ) V(XDUT.vg) V(XDUT.dmem)
.endc
.end
