*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../ciceda/models/ptm_130_ngspice.spi
.include ../../../ciceda/lib/SUN_TR_GF130N.spi
.include ../../../ciceda/lib/SUN_TRIO_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc 1.5
V1 VSTORE VSS dc 0.2 
VSS VSS 0 dc 0

V2 VSTORE VCMP_OUT dc 0

IPB1 VDD VBIAS dc 1u
XMNB0 VBIAS VBIAS VSS VSS NCHCM2

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include comp.cir
XDUT VCMP_OUT VSTORE VRAMP VBIAS VDD VSS COMP

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------

.control
op
* Vds
print v(XDUT.VDIFF1)-v(XDUT.VCURR)
* Vgs
print v(VSTORE)-v(XDUT.VCURR)

* Vgs cm
print v(XDUT.VDIFF1)-v(VDD)

show m.xdut.m1 : vth
show m.xdut.m2 : vth
show m.xdut.m3 : vth
show m.xdut.m4 : vth
.endc
.end
