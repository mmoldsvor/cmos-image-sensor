*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../ciceda/models/ptm_130_ngspice.spi
.include ../../../ciceda/lib/SUN_TR_GF130N.spi
.include ../../../ciceda/lib/SUN_TRIO_GF130N.spi

*----------------------------------------------------------------
* Options
*----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

*----------------------------------------------------------------
* Sources
*----------------------------------------------------------------
VDD VDD VSS dc 1.5
VSS VSS 0 dc 0
VA A VSS PULSE(0, 1.3, 15u, 10n, 10n, 30u, 60u, 0)

*----------------------------------------------------------------
* DUT
*----------------------------------------------------------------
.include xor.cir
X1 A OUT VDD VSS INVERTER

.control
set color0=white
set color1=black
tran 1n 60u
plot V(A) V(OUT)
wrdata ../output/tb_inverter.txt V(A) V(OUT)
.endc
.end