.SUBCKT COMP VIP VIN LATCH OUTP OUTN VDD VSS

M1 COMPOUTP COMPOUTN VDD VDD pmos w=0.5u l=0.5u
M2 COMPOUTN COMPOUTP VDD VDD pmos w=0.5u l=0.5u
M3 COMPOUTP COMPOUTN DIFFP VSS nmos w=0.5u l=0.5u
M4 COMPOUTN COMPOUTP DIFFN VSS nmos w=0.5u l=0.5u

M5 DIFFP VIP DYN VSS nmos w=0.5u l=0.5u
M6 DIFFN VIN DYN VSS nmos w=0.5u l=0.5u

M7 DYN LATCH VSS VSS nmos w=0.5u l=0.5u
M8 DYN LATCH VSS VSS nmos w=0.5u l=0.5u

M9 DIFFP LATCH VDD VDD pmos w=0.5u l=0.5u
M10 COMPOUTP LATCH VDD VDD pmos w=0.5u l=0.5u

M11 DIFFN LATCH VDD VDD pmos w=0.5u l=0.5u
M12 COMPOUTN LATCH VDD VDD pmos w=0.5u l=0.5u

* Inverters
M13 OUTP COMPOUTP VDD VDD pmos w=0.5u l=0.5u
M14 OUTP COMPOUTP VSS VSS nmos w=0.5u l=0.5u
M15 OUTN COMPOUTN VDD VDD pmos w=0.5u l=0.5u
M16 OUTN COMPOUTN VSS VSS nmos w=0.5u l=0.5u

.ENDS