.SUBCKT COMP VCMP_OUT VSTORE VRAMP VBIAS VDD VSS


M3 VDIFF1 VDIFF2 VDD VDD pmos w=0.05u l=0.5u
M4 VDIFF2 VDIFF1 VDD VDD pmos w=0.05u l=0.5u

* Differential pair
M1 VDIFF1 VSTORE VCURR VSS nmos w=1.5u l=0.15u
M2 VDIFF2 VRAMP VCURR VSS nmos w=1.5u l=0.15u

* Current source
XMN3 VCURR VBIAS VSS VSS NCHCM2

* Inverter stage 2
XN5 VINV_OUT VDIFF2 VSS VSS NCH
XP4 VINV_OUT VDIFF2 VDD VDD PCH

* Inverter stage 2
XN6 VCMP_OUT VINV_OUT VSS VSS NCH
XP5 VCMP_OUT VINV_OUT VDD VDD PCH

.ENDS
