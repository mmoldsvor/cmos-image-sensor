.SUBCKT GRAY VDATA0 VDATA1 VDATA2 VDATA3 VDATA4 VDATA5 VDATA6 VDATA7 VOUT0 VOUT1 VOUT2 VOUT3 VOUT4 VOUT5 VOUT6 VOUT7 VDD VSS
    R VDATA7 VOUT7 0
    X1 VDATA7 VDATA6 VOUT6 VDD VSS XOR
    X2 VDATA6 VDATA5 VOUT5 VDD VSS XOR
    X3 VDATA5 VDATA4 VOUT4 VDD VSS XOR
    X4 VDATA4 VDATA3 VOUT3 VDD VSS XOR
    X5 VDATA3 VDATA2 VOUT2 VDD VSS XOR
    X6 VDATA2 VDATA1 VOUT1 VDD VSS XOR
    X7 VDATA1 VDATA0 VOUT0 VDD VSS XOR
.ENDS
