.SUBCKT INVERTER IN OUT VDD VSS
    XP1 OUT IN VDD VDD PCHIO
    XP2 OUT IN VSS VSS NCHIO
.ENDS

.SUBCKT XOR A B OUT VDD VSS
    X1 A A_INV VDD VSS INVERTER
    X2 B B_INV VDD VSS INVERTER

    XP1 LEFT1 A VDD VDD PCHIO
    XP2 OUT B_INV LEFT1 VDD PCHIO
    XN1 OUT A_INV LEFT2 VSS NCHIO
    XN2 LEFT2 B_INV VSS VSS NCHIO

    XP3 RIGHT1 A_INV VDD VDD PCHIO
    XP4 OUT B RIGHT1 VDD PCHIO
    XN3 OUT A RIGHT2 VSS NCHIO
    XN4 RIGHT2 B VSS VSS NCHIO
.ENDS
