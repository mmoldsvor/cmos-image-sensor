.SUBCKT SENSOR VRESET VSTORE ERASE EXPOSE VDD VSS

C1 VSTORE VSS 100f

M1 VRESET ERASE VSTORE VSS nmos w=0.5u l=0.5u

M2 VSTORE EXPOSE VPG VSS nmos w=0.5u l=0.5u

Rphoo VPG VSS 1000Meg
.ENDS