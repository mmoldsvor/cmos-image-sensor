.SUBCKT PIXEL_SENSOR VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

.include sensor.cir
X1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR

.include comp_feedback.cir
X2 VCMP_OUT VSTORE VRAMP VBN1 VDD VSS COMP

.include memory.cir
X3 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY

.ENDS